*** SPICE deck for cell inv{sch} from library Inverter
*** Created on Thu Jun 20, 2024 20:19:54
*** Last revised on Thu Jun 20, 2024 20:49:00
*** Written on Mon Jun 24, 2024 11:56:09 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)

.global gnd vdd

*** TOP LEVEL CELL: inv{sch}
Mnmos@0 out in gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd in out vdd PMOS L=0.4U W=2U

* Spice Code nodes in cell cell 'inv{sch}'
vdd vdd 0 DC 5
vin in 0 DC pwl 10ns 0 20ns 5 50ns 5 60ns 0
cload out 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=8ns targ v(out) val=0.5 fall=1
.measure tran tf trig v(out) val=0.5 rise=1 td=8ns targ v(out) val=4.5 rise=1
.tran 0 0.1us
.include C:\Users\hamza\OneDrive\Documents\electric\C5_models.txt
.END
