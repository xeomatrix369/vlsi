.global gnd vdd

*** TOP LEVEL CELL: nand{sch}
Mnmos@1 net@110 b gnd gnd NMOS L=0.4U W=2U
Mnmos@2 anandb a net@110 gnd NMOS L=0.4U W=2U
Mpmos@0 vdd a anandb vdd PMOS L=0.4U W=2U
Mpmos@1 anandb b vdd vdd PMOS L=0.4U W=2U

* Spice Code nodes in cell cell 'nand{sch}'
vdd vdd 0 DC 5
va a 0 DC pwl 10ns 0 20ns 5 50ns 5 60ns 0 90ns 0 100ns 5 130ns 5 140ns 0 170ns 0 180ns 5
vb b 0 DC pwl 10ns 0 20ns 0 50ns 0 60ns 0 90ns 0 100ns 5 130ns 5 140ns 5 170ns 5 180ns 5
.measure tran tf trig v(anandb) val=4.5 fall=1 td=8ns targ v(out) val=0.5 fall=1
.measure tran tf trig v(anandb) val=0.5 rise=1 td=8ns targ v(out) val=4.5 rise=1
.tran 0 0.2us
.include C:\Users\hamza\OneDrive\Documents\electric\C5_models.txt
.END
