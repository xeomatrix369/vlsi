module buffer (
  input in,
  output out
);

  assign out = in;

endmodule
